netcdf pism_config_override {
variables:
byte pism_overrides;

//beddef
pism_overrides:bed_deformation.lithosphere_flexural_rigidity = 5.0e24;
pism_overrides:bed_deformation.mantle_viscosity = 1.0e21;

//precip
pism_overrides:atmosphere.precip_exponential_factor_for_temperature = .02;

//pdd
pism_overrides:surface.pdd.factor_snow = 3.0e-3;
pism_overrides:surface.pdd.factor_ice = 8.8e-3;
pism_overrides:surface.pdd.std_dev = 5.0;

//sliding
pism_overrides:inverse.ssa.velocity_scale = 100;
pism_overrides:basal_resistance.pseudo_plastic.q = 0.25;
pism_overrides:hydrology.tillwat_decay_rate = 3.16887646154128e-11;
pism_overrides:basal_yield_stress.mohr_coulomb.till_effective_fraction_overburden = 0.02;

//enhancement
pism_overrides:stress_balance.sia.enhancement_factor = 1.0;
pism_overrides:stress_balance.ssa.enhancement_factor = 1.0;

//calving
pism_overrides:calving.eigen_calving.K = 0.0;
pism_overrides:calving.thickness_calving.threshold = 50.0;

//grounding line
pism_overrides:energy.basal_melt.use_grounded_cell_fraction  = "true";
pism_overrides:basal_yield_stress.slippery_grounding_lines = "no";

//topg_to_phi
pism_overrides:basal_yield_stress.mohr_coulomb.topg_to_phi.enabled = "no";
pism_overrides:basal_yield_stress.mohr_coulomb.topg_to_phi.phi_max = 15.0;
pism_overrides:basal_yield_stress.mohr_coulomb.topg_to_phi.phi_min = 5.0;
pism_overrides:basal_yield_stress.mohr_coulomb.topg_to_phi.topg_max = 1000.0;
pism_overrides:basal_yield_stress.mohr_coulomb.topg_to_phi.topg_min = -1000.0;

//pico ocean

//phi optimization

//force_to_thickness

}

//ncgen3 pism_config_override.cdl -o pism_config_override.nc
